LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;
USE work.MyTypes.ALL;

ENTITY testbench IS
    
END testbench;

ARCHITECTURE tb OF testbench IS
	COMPONENT Processor IS
        PORT (
            clk,reset : IN STD_LOGIC
        );
    END COMPONENT;

	signal clk,reset : std_logic;
    
BEGIN

    UUT : Processor PORT MAP(clk,reset);

    PROCESS
    BEGIN
    reset<='1';
    wait for 10 ns;
    reset<='0';
   
    for I in 0 to 40 loop
	    clk <= '0';
        wait for 10 ns;
        clk <= '1';
	    wait for 10 ns;    
    end loop;        
    WAIT;
    END PROCESS;
END tb;